`define CLK_PERIOD 10
`define NUM_BLOCKS 100
`define HRES 320
`define VRES 240
`define HBLOCKS `HRES/16
`define VBLOCKS `VRES/16

`define SIM_BLOCKS 20
