module CoeffTokenLUT02_6 (
                           input [2:0] Bits,
                           output reg [4:0] TotalCoeff, 
                           output reg [1:0] TrailingOnes, 
                           output reg [4:0] NumShift
                           );
always @* begin
  case (Bits)
    3'b110,3'b111 : begin
      TotalCoeff = 5'd3;
      TrailingOnes = 2'd3;
      NumShift = 5'd5;
    end
    3'b101 : begin
      TotalCoeff = 5'd1;
      TrailingOnes = 2'd0;
      NumShift = 5'd6;
    end
    3'b100 : begin
      TotalCoeff = 5'd2;
      TrailingOnes = 2'd1;
      NumShift = 5'd6;
    end
    3'b011 : begin
      TotalCoeff = 5'd4;
      TrailingOnes = 2'd3;
      NumShift = 5'd6;
    end
    default : begin
      TotalCoeff = 'bx;
      TrailingOnes = 'bx;
      NumShift = 'bx;
    end
  endcase
end

endmodule