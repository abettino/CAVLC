`define CLK_PERIOD 10
`define NUM_BLOCKS 100


